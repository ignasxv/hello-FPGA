library verilog;
use verilog.vl_types.all;
entity inv02 is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end inv02;
