library verilog;
use verilog.vl_types.all;
entity test_RTL_multiply is
end test_RTL_multiply;
