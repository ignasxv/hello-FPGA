library verilog;
use verilog.vl_types.all;
entity fake_gnd is
    port(
        Y               : out    vl_logic
    );
end fake_gnd;
