library verilog;
use verilog.vl_types.all;
entity buf02 is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end buf02;
