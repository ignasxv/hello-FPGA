library verilog;
use verilog.vl_types.all;
entity testMultiplier is
end testMultiplier;
