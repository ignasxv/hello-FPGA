library verilog;
use verilog.vl_types.all;
entity testRTL_multiply is
end testRTL_multiply;
