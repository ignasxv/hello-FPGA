// parity adjustemnet test bench

`timescale 1ns/1ps

module test; 
    
endmodule